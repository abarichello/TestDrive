library ieee;
use ieee.std_logic_1164.all;

entity map4 is
	port
	(
		F0, F1, F2, F3, F4, F5, F6, F7, F8, F9, F10, F11, F12, F13, F14, F15: out std_logic_vector(31 downto 0)
	);
end map4;	
	
architecture map4_struct of map4 is
begin
	F0 <=  "00011111111111111111111111000000";
	F1 <=  "00000010000100111111001011000000";
	F2 <=  "00000000000000000000000000000000";
	F3 <=  "00000000000000000000000011000000";
	F4 <=  "00000010000000011100000000000000";
	F5 <=  "00000010000000011100110000000000";
	F6 <=  "00000010000000011100000000000000";
	F7 <=  "00000000000000011100000011000000";
	F8 <=  "00000010000000000100010000000000";
	F9 <=  "00000010000000011100000000000000";
	F10 <= "00000010000000011100000000000000";
	F11 <= "00000010010000000000000000000000";
	F12 <= "00000000000000000000000011000000";
	F13 <= "01001100001111000000100011000000";
	F14 <= "00000000000000011100000011010100";
	F15 <= "00000111111111011100000011000000";
end map4_struct;