library ieee;
use ieee.std_logic_1164.all;

entity map4 is
	port
	(
		F0, F1, F2, F3, F4, F5, F6, F7, F8, F9, F10, F11, F12, F13, F14, F15: out std_logic_vector(31 downto 0)
	);
end map4;	
	
architecture map4_struct of map4 is
begin
	F0 <=  "11011111111111111000111111000110";
	F1 <=  "00000010000111111000101011000000";
	F2 <=  "00000000000011100000000000000000";
	F3 <=  "11100011110000000000111111000001";
	F4 <=  "11110000000000001100000000000001";
	F5 <=  "00000010000000011111110001111100";
	F6 <=  "00000000000000000000000000000000"; --easy lane
	F7 <=  "00000000000010000000000011001100";
	F8 <=  "00000010000000000000010000000011";
	F9 <=  "01110010000000011100000011000011";
	F10 <= "00000000000000011100000011000000";
	F11 <= "10001111010000000000000000000000";
	F12 <= "11000000000100111000000011000000";
	F13 <= "00001100001111111000100111000011";
	F14 <= "10000000000000011100000011010000";
	F15 <= "10011111111111011100111111100000";
end map4_struct;